library ieee;
use ieee.std_logic_1164.all;

package data_types is
    constant screen_w : integer := 640;
    constant screen_h : integer := 480;
    constant img_w : integer := 32;
    constant img_h : integer := 32;
    type IMGTYPE is array (0 to img_w - 1, 0 to img_h - 1) of std_logic_vector (7 downto 0);
    
    constant clr_bmp_w : integer := 88;
    constant clr_bmp_h : integer := 40;
    type CLEAR_BITMAP_TYPE is array (0 to clr_bmp_h - 1, 0 to clr_bmp_w - 1) of std_logic;
    constant clear_bitmap : CLEAR_BITMAP_TYPE := (
        "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "0000000000000000000001111110000011100000000000000000000000000000000000000000000000000000",
        "0000000000000000000011000011000001100000000000000000000000000000000000000000000000000000",
        "0000000000000000000011000011000001100000000000000000000000000000000000000000000000000000",
        "0000000000000000000011000000000001100000011111100001111110001101111100000000000000000000",
        "0000000000000000000011000000000001100000110000110000000011001111000000000000000000000000",
        "0000000000000000000011000000000001100000110000110000000011001110000000000000000000000000",
        "0000000000000000000011000000000001100000110000110001111111001100000000000000000000000000",
        "0000000000000000000011000000000001100000111111110011000011001100000000000000000000000000",
        "0000000000000000000011000000000001100000110000000011000011001100000000000000000000000000",
        "0000000000000000000011000011000001100000110000000011000011001100000000000000000000000000",
        "0000000000000000000011000011000001100000110000110011000011001100000000000000000000000000",
        "0000000000000000000001111110000011110000011111100001111111001100000000000000000000000000",
        "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
        );
end data_types;

package body data_types is

 
end data_types;